module multiplier (
    input A [15:0],
    input B [15:0],
    output result[31:0]
);



endmodule